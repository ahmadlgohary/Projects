library verilog;
use verilog.vl_types.all;
entity controlUnit_vlg_vec_tst is
end controlUnit_vlg_vec_tst;
